------------------------------------------------------------------------------------
---- Company: 
---- Engineer: 
---- 
---- Create Date: 24.12.2024 11:29:47
---- Design Name: 
---- Module Name: unit_operativa - Behavioral
---- Project Name: 
---- Target Devices: 
---- Tool Versions: 
---- Description: 
---- 
---- Dependencies: 
---- 
---- Revision:
---- Revision 0.01 - File Created
---- Additional Comments:
---- 
------------------------------------------------------------------------------------


--library IEEE;
--use IEEE.STD_LOGIC_1164.ALL;

--entity unit_operativa is
----  Port ( );
--end unit_operativa;

--architecture Behavioral of unit_operativa is

--begin


--end Behavioral;
